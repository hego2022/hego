`include "uvm_macros.svh"
`ifndef pkg_svh
`define pkg_svh
package uvm_;
import uvm_pkg::*;
`include "uvm_macros.svh";
endpackage
`endif