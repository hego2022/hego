`include "uvm_macros.svh"
`include "seq item.sv"
import uvm_pkg::*;
class scoreboard extends uvm_subscriber  #(aes_transaction);
   `uvm_component_utils(scoreboard);
   task kat;
bit[127:0] katvk[bit[127:0]];
bit[127:0] katvt [bit[127:0]];
initial
begin
   katvt='{
32'h80000000000000000000000000000000	: 32'h3ad78e726c1ec02b7ebfe92b23d9ec34,
32'hc0000000000000000000000000000000	: 32'haae5939c8efdf2f04e60b9fe7117b2c2,
32'he0000000000000000000000000000000	: 32'hf031d4d74f5dcbf39daaf8ca3af6e527,
32'hf0000000000000000000000000000000	: 32'h96d9fd5cc4f07441727df0f33e401a36,
32'hf8000000000000000000000000000000	: 32'h30ccdb044646d7e1f3ccea3dca08b8c0,
32'hfc000000000000000000000000000000	: 32'h16ae4ce5042a67ee8e177b7c587ecc82,
32'hfe000000000000000000000000000000	: 32'hb6da0bb11a23855d9c5cb1b4c6412e0a,
32'hff000000000000000000000000000000	: 32'hdb4f1aa530967d6732ce4715eb0ee24b,
32'hff800000000000000000000000000000	: 32'ha81738252621dd180a34f3455b4baa2f,
32'hffc00000000000000000000000000000	: 32'h77e2b508db7fd89234caf7939ee5621a,
32'hffe00000000000000000000000000000	: 32'hb8499c251f8442ee13f0933b688fcd19,
32'hfff00000000000000000000000000000	: 32'h965135f8a81f25c9d630b17502f68e53,
32'hfff80000000000000000000000000000	: 32'h8b87145a01ad1c6cede995ea3670454f,
32'hfffc0000000000000000000000000000	: 32'h8eae3b10a0c8ca6d1d3b0fa61e56b0b2,
32'hfffe0000000000000000000000000000	: 32'h64b4d629810fda6bafdf08f3b0d8d2c5,
32'hffff0000000000000000000000000000	: 32'hd7e5dbd3324595f8fdc7d7c571da6c2a,
32'hffff8000000000000000000000000000	: 32'hf3f72375264e167fca9de2c1527d9606,
32'hffffc000000000000000000000000000	: 32'h8ee79dd4f401ff9b7ea945d86666c13b,
32'hffffe000000000000000000000000000	: 32'hdd35cea2799940b40db3f819cb94c08b,
32'hfffff000000000000000000000000000	: 32'h6941cb6b3e08c2b7afa581ebdd607b87,
32'hfffff800000000000000000000000000	: 32'h2c20f439f6bb097b29b8bd6d99aad799,
32'hfffffc00000000000000000000000000	: 32'h625d01f058e565f77ae86378bd2c49b3,
32'hfffffe00000000000000000000000000	: 32'hc0b5fd98190ef45fbb4301438d095950,
32'hffffff00000000000000000000000000	: 32'h13001ff5d99806efd25da34f56be854b,
32'hffffff80000000000000000000000000	: 32'h3b594c60f5c8277a5113677f94208d82,
32'hffffffc0000000000000000000000000	: 32'he9c0fc1818e4aa46bd2e39d638f89e05,
32'hffffffe0000000000000000000000000	: 32'hf8023ee9c3fdc45a019b4e985c7e1a54,
32'hfffffff0000000000000000000000000	: 32'h35f40182ab4662f3023baec1ee796b57,
32'hfffffff8000000000000000000000000	: 32'h3aebbad7303649b4194a6945c6cc3694,
32'hfffffffc000000000000000000000000	: 32'ha2124bea53ec2834279bed7f7eb0f938,
32'hfffffffe000000000000000000000000	: 32'hb9fb4399fa4facc7309e14ec98360b0a,
32'hffffffff000000000000000000000000	: 32'hc26277437420c5d634f715aea81a9132,
32'hffffffff800000000000000000000000	: 32'h171a0e1b2dd424f0e089af2c4c10f32f,
32'hffffffffc00000000000000000000000	: 32'h7cadbe402d1b208fe735edce00aee7ce,
32'hffffffffe00000000000000000000000	: 32'h43b02ff929a1485af6f5c6d6558baa0f,
32'hfffffffff00000000000000000000000	: 32'h092faacc9bf43508bf8fa8613ca75dea,
32'hfffffffff80000000000000000000000	: 32'hcb2bf8280f3f9742c7ed513fe802629c,
32'hfffffffffc0000000000000000000000	: 32'h215a41ee442fa992a6e323986ded3f68,
32'hfffffffffe0000000000000000000000	: 32'hf21e99cf4f0f77cea836e11a2fe75fb1,
32'hffffffffff0000000000000000000000	: 32'h95e3a0ca9079e646331df8b4e70d2cd6,
32'hffffffffff8000000000000000000000	: 32'h4afe7f120ce7613f74fc12a01a828073,
32'hffffffffffc000000000000000000000	: 32'h827f000e75e2c8b9d479beed913fe678,
32'hffffffffffe000000000000000000000	: 32'h35830c8e7aaefe2d30310ef381cbf691,
32'hfffffffffff000000000000000000000	: 32'h191aa0f2c8570144f38657ea4085ebe5,
32'hfffffffffff800000000000000000000	: 32'h85062c2c909f15d9269b6c18ce99c4f0,
32'hfffffffffffc00000000000000000000	: 32'h678034dc9e41b5a560ed239eeab1bc78,
32'hfffffffffffe00000000000000000000	: 32'hc2f93a4ce5ab6d5d56f1b93cf19911c1,
32'hffffffffffff00000000000000000000	: 32'h1c3112bcb0c1dcc749d799743691bf82,
32'hffffffffffff80000000000000000000	: 32'h00c55bd75c7f9c881989d3ec1911c0d4,
32'hffffffffffffc0000000000000000000	: 32'hea2e6b5ef182b7dff3629abd6a12045f,
32'hffffffffffffe0000000000000000000	: 32'h22322327e01780b17397f24087f8cc6f,
32'hfffffffffffff0000000000000000000	: 32'hc9cacb5cd11692c373b2411768149ee7,
32'hfffffffffffff8000000000000000000	: 32'ha18e3dbbca577860dab6b80da3139256,
32'hfffffffffffffc000000000000000000	: 32'h79b61c37bf328ecca8d743265a3d425c,
32'hfffffffffffffe000000000000000000	: 32'hd2d99c6bcc1f06fda8e27e8ae3f1ccc7,
32'hffffffffffffff000000000000000000	: 32'h1bfd4b91c701fd6b61b7f997829d663b,
32'hffffffffffffff800000000000000000	: 32'h11005d52f25f16bdc9545a876a63490a,
32'hffffffffffffffc00000000000000000	: 32'h3a4d354f02bb5a5e47d39666867f246a,
32'hffffffffffffffe00000000000000000	: 32'hd451b8d6e1e1a0ebb155fbbf6e7b7dc3,
32'hfffffffffffffff00000000000000000	: 32'h6898d4f42fa7ba6a10ac05e87b9f2080,
32'hfffffffffffffff80000000000000000	: 32'hb611295e739ca7d9b50f8e4c0e754a3f,
32'hfffffffffffffffc0000000000000000	: 32'h7d33fc7d8abe3ca1936759f8f5deaf20,
32'hfffffffffffffffe0000000000000000	: 32'h3b5e0f566dc96c298f0c12637539b25c,
32'hffffffffffffffff0000000000000000	: 32'hf807c3e7985fe0f5a50e2cdb25c5109e,
32'hffffffffffffffff8000000000000000	: 32'h41f992a856fb278b389a62f5d274d7e9,
32'hffffffffffffffffc000000000000000	: 32'h10d3ed7a6fe15ab4d91acbc7d0767ab1,
32'hffffffffffffffffe000000000000000	: 32'h21feecd45b2e675973ac33bf0c5424fc,
32'hfffffffffffffffff000000000000000	: 32'h1480cb3955ba62d09eea668f7c708817,
32'hfffffffffffffffff800000000000000	: 32'h66404033d6b72b609354d5496e7eb511,
32'hfffffffffffffffffc00000000000000	: 32'h1c317a220a7d700da2b1e075b00266e1,
32'hfffffffffffffffffe00000000000000	: 32'hab3b89542233f1271bf8fd0c0f403545,
32'hffffffffffffffffff00000000000000	: 32'hd93eae966fac46dca927d6b114fa3f9e,
32'hffffffffffffffffff80000000000000	: 32'h1bdec521316503d9d5ee65df3ea94ddf,
32'hffffffffffffffffffc0000000000000	: 32'heef456431dea8b4acf83bdae3717f75f,
32'hffffffffffffffffffe0000000000000	: 32'h06f2519a2fafaa596bfef5cfa15c21b9,
32'hfffffffffffffffffff0000000000000	: 32'h251a7eac7e2fe809e4aa8d0d7012531a,
32'hfffffffffffffffffff8000000000000	: 32'h3bffc16e4c49b268a20f8d96a60b4058,
32'hfffffffffffffffffffc000000000000	: 32'he886f9281999c5bb3b3e8862e2f7c988,
32'hfffffffffffffffffffe000000000000	: 32'h563bf90d61beef39f48dd625fcef1361,
32'hffffffffffffffffffff000000000000	: 32'h4d37c850644563c69fd0acd9a049325b,
32'hffffffffffffffffffff800000000000	: 32'hb87c921b91829ef3b13ca541ee1130a6,
32'hffffffffffffffffffffc00000000000	: 32'h2e65eb6b6ea383e109accce8326b0393,
32'hffffffffffffffffffffe00000000000	: 32'h9ca547f7439edc3e255c0f4d49aa8990,
32'hfffffffffffffffffffff00000000000	: 32'ha5e652614c9300f37816b1f9fd0c87f9,
32'hfffffffffffffffffffff80000000000	: 32'h14954f0b4697776f44494fe458d814ed,
32'hfffffffffffffffffffffc0000000000	: 32'h7c8d9ab6c2761723fe42f8bb506cbcf7,
32'hfffffffffffffffffffffe0000000000	: 32'hdb7e1932679fdd99742aab04aa0d5a80,
32'hffffffffffffffffffffff0000000000	: 32'h4c6a1c83e568cd10f27c2d73ded19c28,
32'hffffffffffffffffffffff8000000000	: 32'h90ecbe6177e674c98de412413f7ac915,
32'hffffffffffffffffffffffc000000000	: 32'h90684a2ac55fe1ec2b8ebd5622520b73,
32'hffffffffffffffffffffffe000000000	: 32'h7472f9a7988607ca79707795991035e6,
32'hfffffffffffffffffffffff000000000	: 32'h56aff089878bf3352f8df172a3ae47d8,
32'hfffffffffffffffffffffff800000000	: 32'h65c0526cbe40161b8019a2a3171abd23,
32'hfffffffffffffffffffffffc00000000	: 32'h377be0be33b4e3e310b4aabda173f84f,
32'hfffffffffffffffffffffffe00000000	: 32'h9402e9aa6f69de6504da8d20c4fcaa2f,
32'hffffffffffffffffffffffff00000000	: 32'h123c1f4af313ad8c2ce648b2e71fb6e1,
32'hffffffffffffffffffffffff80000000	: 32'h1ffc626d30203dcdb0019fb80f726cf4,
32'hffffffffffffffffffffffffc0000000	: 32'h76da1fbe3a50728c50fd2e621b5ad885,
32'hffffffffffffffffffffffffe0000000	: 32'h082eb8be35f442fb52668e16a591d1d6,
32'hfffffffffffffffffffffffff0000000	: 32'he656f9ecf5fe27ec3e4a73d00c282fb3,
32'hfffffffffffffffffffffffff8000000	: 32'h2ca8209d63274cd9a29bb74bcd77683a,
32'hfffffffffffffffffffffffffc000000	: 32'h79bf5dce14bb7dd73a8e3611de7ce026,
32'hfffffffffffffffffffffffffe000000	: 32'h3c849939a5d29399f344c4a0eca8a576,
32'hffffffffffffffffffffffffff000000	: 32'hed3c0a94d59bece98835da7aa4f07ca2,
32'hffffffffffffffffffffffffff800000	: 32'h63919ed4ce10196438b6ad09d99cd795,
32'hffffffffffffffffffffffffffc00000	: 32'h7678f3a833f19fea95f3c6029e2bc610,
32'hffffffffffffffffffffffffffe00000	: 32'h3aa426831067d36b92be7c5f81c13c56,
32'hfffffffffffffffffffffffffff00000	: 32'h9272e2d2cdd11050998c845077a30ea0,
32'hfffffffffffffffffffffffffff80000	: 32'h088c4b53f5ec0ff814c19adae7f6246c,
32'hfffffffffffffffffffffffffffc0000	: 32'h4010a5e401fdf0a0354ddbcc0d012b17,
32'hfffffffffffffffffffffffffffe0000	: 32'ha87a385736c0a6189bd6589bd8445a93,
32'hffffffffffffffffffffffffffff0000	: 32'h545f2b83d9616dccf60fa9830e9cd287,
32'hffffffffffffffffffffffffffff8000	: 32'h4b706f7f92406352394037a6d4f4688d,
32'hffffffffffffffffffffffffffffc000	: 32'hb7972b3941c44b90afa7b264bfba7387,
32'hffffffffffffffffffffffffffffe000	: 32'h6f45732cf10881546f0fd23896d2bb60,
32'hfffffffffffffffffffffffffffff000	: 32'h2e3579ca15af27f64b3c955a5bfc30ba,
32'hfffffffffffffffffffffffffffff800	: 32'h34a2c5a91ae2aec99b7d1b5fa6780447,
32'hfffffffffffffffffffffffffffffc00	: 32'ha4d6616bd04f87335b0e53351227a9ee,
32'hfffffffffffffffffffffffffffffe00	: 32'h7f692b03945867d16179a8cefc83ea3f,
32'hffffffffffffffffffffffffffffff00	: 32'h3bd141ee84a0e6414a26e7a4f281f8a2,
32'hffffffffffffffffffffffffffffff80	: 32'hd1788f572d98b2b16ec5d5f3922b99bc,
32'hffffffffffffffffffffffffffffffc0	: 32'h0833ff6f61d98a57b288e8c3586b85a6,
32'hffffffffffffffffffffffffffffffe0	: 32'h8568261797de176bf0b43becc6285afb,
32'hfffffffffffffffffffffffffffffff0	: 32'hf9b0fda0c4a898f5b9e6f661c4ce4d07,
32'hfffffffffffffffffffffffffffffff8	: 32'h8ade895913685c67c5269f8aae42983e,
32'hfffffffffffffffffffffffffffffffc	: 32'h39bde67d5c8ed8a8b1c37eb8fa9f5ac0,
32'hfffffffffffffffffffffffffffffffe	: 32'h5c005e72c1418c44f569f2ea33ba54f3,
32'hffffffffffffffffffffffffffffffff	: 32'h3f5b8cc9ea855a0afa7347d23e8d664e
};
   katvk='{
32'h80000000000000000000000000000000	: 32'h0edd33d3c621e546455bd8ba1418bec8,
32'hc0000000000000000000000000000000	: 32'h4bc3f883450c113c64ca42e1112a9e87,
32'he0000000000000000000000000000000	: 32'h72a1da770f5d7ac4c9ef94d822affd97,
32'hf0000000000000000000000000000000	: 32'h970014d634e2b7650777e8e84d03ccd8,
32'hf8000000000000000000000000000000	: 32'hf17e79aed0db7e279e955b5f493875a7,
32'hfc000000000000000000000000000000	: 32'h9ed5a75136a940d0963da379db4af26a,
32'hfe000000000000000000000000000000	: 32'hc4295f83465c7755e8fa364bac6a7ea5,
32'hff000000000000000000000000000000	: 32'hb1d758256b28fd850ad4944208cf1155,
32'hff800000000000000000000000000000	: 32'h42ffb34c743de4d88ca38011c990890b,
32'hffc00000000000000000000000000000	: 32'h9958f0ecea8b2172c0c1995f9182c0f3,
32'hffe00000000000000000000000000000	: 32'h956d7798fac20f82a8823f984d06f7f5,
32'hfff00000000000000000000000000000	: 32'ha01bf44f2d16be928ca44aaf7b9b106b,
32'hfff80000000000000000000000000000	: 32'hb5f1a33e50d40d103764c76bd4c6b6f8,
32'hfffc0000000000000000000000000000	: 32'h2637050c9fc0d4817e2d69de878aee8d,
32'hfffe0000000000000000000000000000	: 32'h113ecbe4a453269a0dd26069467fb5b5,
32'hffff0000000000000000000000000000	: 32'h97d0754fe68f11b9e375d070a608c884,
32'hffff8000000000000000000000000000	: 32'hc6a0b3e998d05068a5399778405200b4,
32'hffffc000000000000000000000000000	: 32'hdf556a33438db87bc41b1752c55e5e49,
32'hffffe000000000000000000000000000	: 32'h90fb128d3a1af6e548521bb962bf1f05,
32'hfffff000000000000000000000000000	: 32'h26298e9c1db517c215fadfb7d2a8d691,
32'hfffff800000000000000000000000000	: 32'ha6cb761d61f8292d0df393a279ad0380,
32'hfffffc00000000000000000000000000	: 32'h12acd89b13cd5f8726e34d44fd486108,
32'hfffffe00000000000000000000000000	: 32'h95b1703fc57ba09fe0c3580febdd7ed4,
32'hffffff00000000000000000000000000	: 32'hde11722d893e9f9121c381becc1da59a,
32'hffffff80000000000000000000000000	: 32'h6d114ccb27bf391012e8974c546d9bf2,
32'hffffffc0000000000000000000000000	: 32'h5ce37e17eb4646ecfac29b9cc38d9340,
32'hffffffe0000000000000000000000000	: 32'h18c1b6e2157122056d0243d8a165cddb,
32'hfffffff0000000000000000000000000	: 32'h99693e6a59d1366c74d823562d7e1431,
32'hfffffff8000000000000000000000000	: 32'h6c7c64dc84a8bba758ed17eb025a57e3,
32'hfffffffc000000000000000000000000	: 32'he17bc79f30eaab2fac2cbbe3458d687a,
32'hfffffffe000000000000000000000000	: 32'h1114bc2028009b923f0b01915ce5e7c4,
32'hffffffff000000000000000000000000	: 32'h9c28524a16a1e1c1452971caa8d13476,
32'hffffffff800000000000000000000000	: 32'hed62e16363638360fdd6ad62112794f0,
32'hffffffffc00000000000000000000000	: 32'h5a8688f0b2a2c16224c161658ffd4044,
32'hffffffffe00000000000000000000000	: 32'h23f710842b9bb9c32f26648c786807ca,
32'hfffffffff00000000000000000000000	: 32'h44a98bf11e163f632c47ec6a49683a89,
32'hfffffffff80000000000000000000000	: 32'h0f18aff94274696d9b61848bd50ac5e5,
32'hfffffffffc0000000000000000000000	: 32'h82408571c3e2424540207f833b6dda69,
32'hfffffffffe0000000000000000000000	: 32'h303ff996947f0c7d1f43c8f3027b9b75,
32'hffffffffff0000000000000000000000	: 32'h7df4daf4ad29a3615a9b6ece5c99518a,
32'hffffffffff8000000000000000000000	: 32'hc72954a48d0774db0b4971c526260415,
32'hffffffffffc000000000000000000000	: 32'h1df9b76112dc6531e07d2cfda04411f0,
32'hffffffffffe000000000000000000000	: 32'h8e4d8e699119e1fc87545a647fb1d34f,
32'hfffffffffff000000000000000000000	: 32'he6c4807ae11f36f091c57d9fb68548d1,
32'hfffffffffff800000000000000000000	: 32'h8ebf73aad49c82007f77a5c1ccec6ab4,
32'hfffffffffffc00000000000000000000	: 32'h4fb288cc2040049001d2c7585ad123fc,
32'hfffffffffffe00000000000000000000	: 32'h04497110efb9dceb13e2b13fb4465564,
32'hffffffffffff00000000000000000000	: 32'h75550e6cb5a88e49634c9ab69eda0430,
32'hffffffffffff80000000000000000000	: 32'hb6768473ce9843ea66a81405dd50b345,
32'hffffffffffffc0000000000000000000	: 32'hcb2f430383f9084e03a653571e065de6,
32'hffffffffffffe0000000000000000000	: 32'hff4e66c07bae3e79fb7d210847a3b0ba,
32'hfffffffffffff0000000000000000000	: 32'h7b90785125505fad59b13c186dd66ce3,
32'hfffffffffffff8000000000000000000	: 32'h8b527a6aebdaec9eaef8eda2cb7783e5,
32'hfffffffffffffc000000000000000000	: 32'h43fdaf53ebbc9880c228617d6a9b548b,
32'hfffffffffffffe000000000000000000	: 32'h53786104b9744b98f052c46f1c850d0b,
32'hffffffffffffff000000000000000000	: 32'hb5ab3013dd1e61df06cbaf34ca2aee78,
32'hffffffffffffff800000000000000000	: 32'h7470469be9723030fdcc73a8cd4fbb10,
32'hffffffffffffffc00000000000000000	: 32'ha35a63f5343ebe9ef8167bcb48ad122e,
32'hffffffffffffffe00000000000000000	: 32'hfd8687f0757a210e9fdf181204c30863,
32'hfffffffffffffff00000000000000000	: 32'h7a181e84bd5457d26a88fbae96018fb0,
32'hfffffffffffffff80000000000000000	: 32'h653317b9362b6f9b9e1a580e68d494b5,
32'hfffffffffffffffc0000000000000000	: 32'h995c9dc0b689f03c45867b5faa5c18d1,
32'hfffffffffffffffe0000000000000000	: 32'h77a4d96d56dda398b9aabecfc75729fd,
32'hffffffffffffffff0000000000000000	: 32'h84be19e053635f09f2665e7bae85b42d,
32'hffffffffffffffff8000000000000000	: 32'h32cd652842926aea4aa6137bb2be2b5e,
32'hffffffffffffffffc000000000000000	: 32'h493d4a4f38ebb337d10aa84e9171a554,
32'hffffffffffffffffe000000000000000	: 32'hd9bff7ff454b0ec5a4a2a69566e2cb84,
32'hfffffffffffffffff000000000000000	: 32'h3535d565ace3f31eb249ba2cc6765d7a,
32'hfffffffffffffffff800000000000000	: 32'hf60e91fc3269eecf3231c6e9945697c6,
32'hfffffffffffffffffc00000000000000	: 32'hab69cfadf51f8e604d9cc37182f6635a,
32'hfffffffffffffffffe00000000000000	: 32'h7866373f24a0b6ed56e0d96fcdafb877,
32'hffffffffffffffffff00000000000000	: 32'h1ea448c2aac954f5d812e9d78494446a,
32'hffffffffffffffffff80000000000000	: 32'hacc5599dd8ac02239a0fef4a36dd1668,
32'hffffffffffffffffffc0000000000000	: 32'hd8764468bb103828cf7e1473ce895073,
32'hffffffffffffffffffe0000000000000	: 32'h1b0d02893683b9f180458e4aa6b73982,
32'hfffffffffffffffffff0000000000000	: 32'h96d9b017d302df410a937dcdb8bb6e43,
32'hfffffffffffffffffff8000000000000	: 32'hef1623cc44313cff440b1594a7e21cc6,
32'hfffffffffffffffffffc000000000000	: 32'h284ca2fa35807b8b0ae4d19e11d7dbd7,
32'hfffffffffffffffffffe000000000000	: 32'hf2e976875755f9401d54f36e2a23a594,
32'hffffffffffffffffffff000000000000	: 32'hec198a18e10e532403b7e20887c8dd80,
32'hffffffffffffffffffff800000000000	: 32'h545d50ebd919e4a6949d96ad47e46a80,
32'hffffffffffffffffffffc00000000000	: 32'hdbdfb527060e0a71009c7bb0c68f1d44,
32'hffffffffffffffffffffe00000000000	: 32'h9cfa1322ea33da2173a024f2ff0d896d,
32'hfffffffffffffffffffff00000000000	: 32'h8785b1a75b0f3bd958dcd0e29318c521,
32'hfffffffffffffffffffff80000000000	: 32'h38f67b9e98e4a97b6df030a9fcdd0104,
32'hfffffffffffffffffffffc0000000000	: 32'h192afffb2c880e82b05926d0fc6c448b,
32'hfffffffffffffffffffffe0000000000	: 32'h6a7980ce7b105cf530952d74daaf798c,
32'hffffffffffffffffffffff0000000000	: 32'hea3695e1351b9d6858bd958cf513ef6c,
32'hffffffffffffffffffffff8000000000	: 32'h6da0490ba0ba0343b935681d2cce5ba1,
32'hffffffffffffffffffffffc000000000	: 32'hf0ea23af08534011c60009ab29ada2f1,
32'hffffffffffffffffffffffe000000000	: 32'hff13806cf19cc38721554d7c0fcdcd4b,
32'hfffffffffffffffffffffff000000000	: 32'h6838af1f4f69bae9d85dd188dcdf0688,
32'hfffffffffffffffffffffff800000000	: 32'h36cf44c92d550bfb1ed28ef583ddf5d7,
32'hfffffffffffffffffffffffc00000000	: 32'hd06e3195b5376f109d5c4ec6c5d62ced,
32'hfffffffffffffffffffffffe00000000	: 32'hc440de014d3d610707279b13242a5c36,
32'hffffffffffffffffffffffff00000000	: 32'hf0c5c6ffa5e0bd3a94c88f6b6f7c16b9,
32'hffffffffffffffffffffffff80000000	: 32'h3e40c3901cd7effc22bffc35dee0b4d9,
32'hffffffffffffffffffffffffc0000000	: 32'hb63305c72bedfab97382c406d0c49bc6,
32'hffffffffffffffffffffffffe0000000	: 32'h36bbaab22a6bd4925a99a2b408d2dbae,
32'hfffffffffffffffffffffffff0000000	: 32'h307c5b8fcd0533ab98bc51e27a6ce461,
32'hfffffffffffffffffffffffff8000000	: 32'h829c04ff4c07513c0b3ef05c03e337b5,
32'hfffffffffffffffffffffffffc000000	: 32'hf17af0e895dda5eb98efc68066e84c54,
32'hfffffffffffffffffffffffffe000000	: 32'h277167f3812afff1ffacb4a934379fc3,
32'hffffffffffffffffffffffffff000000	: 32'h2cb1dc3a9c72972e425ae2ef3eb597cd,
32'hffffffffffffffffffffffffff800000	: 32'h36aeaa3a213e968d4b5b679d3a2c97fe,
32'hffffffffffffffffffffffffffc00000	: 32'h9241daca4fdd034a82372db50e1a0f3f,
32'hffffffffffffffffffffffffffe00000	: 32'hc14574d9cd00cf2b5a7f77e53cd57885,
32'hfffffffffffffffffffffffffff00000	: 32'h793de39236570aba83ab9b737cb521c9,
32'hfffffffffffffffffffffffffff80000	: 32'h16591c0f27d60e29b85a96c33861a7ef,
32'hfffffffffffffffffffffffffffc0000	: 32'h44fb5c4d4f5cb79be5c174a3b1c97348,
32'hfffffffffffffffffffffffffffe0000	: 32'h674d2b61633d162be59dde04222f4740,
32'hffffffffffffffffffffffffffff0000	: 32'hb4750ff263a65e1f9e924ccfd98f3e37,
32'hffffffffffffffffffffffffffff8000	: 32'h62d0662d6eaeddedebae7f7ea3a4f6b6,
32'hffffffffffffffffffffffffffffc000	: 32'h70c46bb30692be657f7eaa93ebad9897,
32'hffffffffffffffffffffffffffffe000	: 32'h323994cfb9da285a5d9642e1759b224a,
32'hfffffffffffffffffffffffffffff000	: 32'h1dbf57877b7b17385c85d0b54851e371,
32'hfffffffffffffffffffffffffffff800	: 32'hdfa5c097cdc1532ac071d57b1d28d1bd,
32'hfffffffffffffffffffffffffffffc00	: 32'h3a0c53fa37311fc10bd2a9981f513174,
32'hfffffffffffffffffffffffffffffe00	: 32'hba4f970c0a25c41814bdae2e506be3b4,
32'hffffffffffffffffffffffffffffff00	: 32'h2dce3acb727cd13ccd76d425ea56e4f6,
32'hffffffffffffffffffffffffffffff80	: 32'h5160474d504b9b3eefb68d35f245f4b3,
32'hffffffffffffffffffffffffffffffc0	: 32'h41a8a947766635dec37553d9a6c0cbb7,
32'hffffffffffffffffffffffffffffffe0	: 32'h25d6cfe6881f2bf497dd14cd4ddf445b,
32'hfffffffffffffffffffffffffffffff0	: 32'h41c78c135ed9e98c096640647265da1e,
32'hfffffffffffffffffffffffffffffff8	: 32'h5a4d404d8917e353e92a21072c3b2305,
32'hfffffffffffffffffffffffffffffffc	: 32'h02bc96846b3fdc71643f384cd3cc3eaf,
32'hfffffffffffffffffffffffffffffffe	: 32'h9ba4a9143f4e5d4048521c4f8877d88e,
32'hffffffffffffffffffffffffffffffff	: 32'ha1f6258c877d5fcd8964484538bfc92c
};
end
endtask
        uvm_analysis_export #(aes_transaction) export_before;
	uvm_analysis_export #(aes_transaction) export_after;

	uvm_tlm_analysis_fifo #(aes_transaction) before_fifo;
	uvm_tlm_analysis_fifo #(aes_transaction) after_fifo;

   
   function new (string name, uvm_component parent);
      super.new(name, parent);
   endfunction : new

   function void build_phase(uvm_phase phase);
      fifo = new ("fifo", this);
   endfunction : build_phase

    function void connect_phase(uvm_phase phase);
	export_before.connect(before_fifo.analysis_export);
	export_after.connect(after_fifo.analysis_export);
    endfunction:connect_phase

   parameter N=99;
   bit[127:0] ct_mc[99:0],pt_mc[99:0],k_mc[99:0];
   bit[127:0] ct_mm[9:0],pt_mm[9:0],k_mm[9:0];
   //function to scan the test vectors
   function read_file(string location,bit[127:0] ct[N:0],pt[N:0],k[N:0]);
      int c,fd,m;
      fd = $fopen(location,"r");
       while(!$feof(fd))
         begin
          m=$fscanf(fd,"COUNT = %d\n",c);
          m=$fscanf(fd,"KEY = %h\n",k[c]);
          m=$fscanf(fd,"PLAINTEXT = %h\n",pt[c]);
          m=$fscanf(fd,"CIPHERTEXT = %h\n\n",ct[c]);
         $display(" %d\n %h\n %h\n %h",c,k[c],pt[c],ct[c]);
         end
   endfunction
//function to extract the result from the test vectors
function  predict_result(aes_transaction cmd);
   bit[127:0] ct_mc[99:0],pt_mc[99:0],k_mc[99:0];
      bit[127:0] predicted;
   if(cmd.opcode_i==AESENCFULL)
    begin
    if(cmd.aes_128 key_i==0)
    predicted=katvt[cmd.aes_128 plain_text_i];
	 else if(cmd.aes_128 plain_text_i==0)
	 predicted=katvk[cmd.aes_128 key_i];
	 else
	 begin
	 read_file("ECBMCT128.txt",ct_mc,pt_mc,k_mc);
	 if(pt_mc.exists(cmd.aes_128 plain_text_i)&&k_mc.exists(cmd.aes_128 key_i))
	 predicted=ct_mc[pt_mc.find_index with (item=aes_128 plain_text_i0];
	 else
	  // where i should put the mmt 
	 end
   end 

   return predicted;
compare();
endfunction : predict_result
 
  virtual function void compare();
		if(aes_transaction == predicted) begin
			`uvm_info("compare", {"Test: OK!"}, UVM_LOW);
		end else begin
			`uvm_error("compare", {"Test: Fail!"}, UVM_LOW);
		end
	endfunction: compare



  endclass : scoreboard

