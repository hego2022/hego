`include "uvm_macros.svh"
`ifndef env_svh
`define env_svh
import uvm_pkg::*;
class env extends uvm_env ;
`uvm_component_utils(env);
endclass
`endif